library verilog;
use verilog.vl_types.all;
entity risc16ba_sv_unit is
end risc16ba_sv_unit;
