library verilog;
use verilog.vl_types.all;
entity sim_risc16ba is
end sim_risc16ba;
